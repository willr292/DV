library verilog;
use verilog.vl_types.all;
entity example_calc1_tb is
end example_calc1_tb;
